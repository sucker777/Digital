library verilog;
use verilog.vl_types.all;
entity Poker_vlg_vec_tst is
end Poker_vlg_vec_tst;
