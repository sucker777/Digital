library verilog;
use verilog.vl_types.all;
entity Poker_Controller_vlg_vec_tst is
end Poker_Controller_vlg_vec_tst;
